module hello_world; 
initial begin
  $display("Hello world!");
  #20 $finish;
end
  
endmodule
